// Copyright 2016 Tudor Timisescu (verificationgentleman.com)
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//     http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.


package reflection;
  import vpi::*;

  `include "reflection_types.svh"

  `include "reflection_rf_value.svh"
  `include "reflection_rf_object_instance.svh"
  `include "reflection_rf_variable.svh"
  `include "reflection_rf_io_declaration.svh"
  `include "reflection_rf_method.svh"
  `include "reflection_rf_task.svh"
  `include "reflection_rf_function.svh"
  `include "reflection_rf_class.svh"
  `include "reflection_rf_package.svh"
  `include "reflection_rf_manager.svh"
endpackage
